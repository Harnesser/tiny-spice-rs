Full-Wave Rectifier with parameterised subcircuits

* 3 instances of a diode bridge + RC load
* cap load in each instances parameterised and overriden from
*   the toplevel

V1 vstack1 gnd     SIN(0 5 1e3) ; input voltage
V2 vstack2 vstack1 SIN(0 2 2e3)
V3 IN_p vstack2    SIN(0 1 3e3)

* full-wave rectifier
.subckt bridge bp bn ba bb

  D1 bp ba
  D2 bb bp
  D3 bn ba
  D4 bb bn

  * Small caps across the diodes to prevent time-step-too-small
  CD1 bp ba 12pF
  CD2 bb bp 12pF
  CD3 bn ba 12pF
  CD4 bb bn 12pF

.ends

.subckt system sinp sinn soutp soutn cval=10uF
  Xbridge sinp sinn midnode soutn bridge
  Rd midnode soutp 1
  Xload soutp soutn r_load cval={cval}
.ends

* Load
.subckt r_load in1 in2 cval=1nF
* Split R so we have internal nodes
  Rl1 in1 la 200
  Rl2 la lb 300
  Rl3 lb lc 400
  Rl4 lc in2 100
  Cload in1 in2 {cval}
.ends

Xsystem1 IN_p gnd vp1 vn1 system cval=1uF
Xsystem2 IN_p gnd vp2 vn2 system cval=10uF
Xsystem3 IN_p gnd vp3 vn3 system cval=100uF

.control
*  option reltol = 0.001
*  option abstol = 1e-12

  tran 100ns 5ms
  option ; ngspice only shows new values after analysis

  plot v(IN_p) v(vp1,vn1) v(vp2,vn2) v(vp3,vn3); (ngspice)
.endc
